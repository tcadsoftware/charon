THIS CIRCUIT IS A MOS LEVEL 1 MODEL CMOS INVERTER AND USES A PARASITIC RESISTOR

VDDdev VDD   0 5V
RIN     IN   1 1K
VIN1     1   0 4.0V

***********************
* one contact version *
***********************
*R1     VOUT  0 10k
***********************
vcr    VOUT  0 0.5
***********************

***********************
* two contact version *
***********************
*R1      VOUT VO 5
*R2       VOO  0 5
***********************
*vcl     VOO   0 0.5
*vcr      VO   0 0.5
***********************

C2    VOUT   0 0.1p
MN1   VOUT  IN   0   0 CD4012_NMOS L=5u W=175u
MP1   VOUT  IN VDD VDD CD4012_PMOS L=5u W=270u

.MODEL cd4012_pmos PMOS
.MODEL cd4012_nmos NMOS

.DC VIN1 0 5 0.5
*.PRINT DC V(vout) v(in) i(R1)
.PRINT DC V(vout) v(in)

.options nonlin nox=1
.options device debuglevel=-100
.END