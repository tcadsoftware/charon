Resistor Circuit Netlist - lower level.
********************************************************************************
R1          1 2 30
VL          1 0 1.0
vconnectR   2 0 0.4
.DC VL 5 5 0
.options nonlin nox=1 
.options device debuglevel=-100
.print dc I(VL) I(vconnectR)
.END