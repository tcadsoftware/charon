Resistor Circuit Netlist - lower level.
********************************************************************************
R1          1 2 3
vconnectL   2 0 1.0
vconnectR   3 0 3.0
R2          3 0 5
vswept      1 0 5.0
.DC vswept 5 5 0
.options nonlin nox=1 
.options device debuglevel=-100
.END

